`include "defines.sv"
`include "multiplexer.sv"
`include "SHFL.sv"
`include "ALU.sv"
