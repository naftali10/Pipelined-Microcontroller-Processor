`define ALU_OP_AMT 8
