`include "defines.sv"		// has to be first
`include "multiplexer.sv"
`include "SHFL.sv"
`include "ALU.sv"
`include "RF.sv"
`include "controller.sv"
